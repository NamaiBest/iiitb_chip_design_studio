/home/vlsiuser/Desktop/team_friday/Cadence_design_database_45nm/Cadence_design_database_45nm/lef/gsclib045_macro.lef