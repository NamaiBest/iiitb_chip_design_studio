/home/vlsiuser21/Downloads/files_rtl3gds/Cadence_design_database_45nm/Cadence_design_database_45nm/lef/gsclib045_macro.lef