/home/vlsiuser/Desktop/team_friday_week2/Cadence_design_database_45nm/Cadence_design_database_45nm/lef/gsclib045_macro.lef